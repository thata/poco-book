module adder(
    input a, b,
    output s);

    assign s = a + b;
endmodule
